LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity process_unit is
    port (  clk : in std_logic;
            key : in std_logic_vector(1 downto 0);
         );
end entity;

architecture rtl of process_unit is
begin
end architecture;
